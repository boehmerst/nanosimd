library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.nanosimd_pkg.all;
use work.func_pkg.all;

entity iexecute is
end entity iexecute;

architecture rtl of iexecute is
begin
end architecture rtl;

